module steering(left, right, walk, sensors);
    output 	left, right, walk;
    input [4:0] 	sensors;
   

endmodule // steering
